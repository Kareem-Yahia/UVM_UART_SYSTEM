 class sys_scoreboard_3 extends uvm_component;
     `uvm_component_utils(sys_scoreboard_3)
 
     function new (string name = "sys_scoreboard_3", uvm_component parent = null);
         super.new(name, parent);
     endfunction
 
 endclass