 
class sys_scoreboard_1 extends uvm_scoreboard;
     `uvm_component_utils(sys_scoreboard_1)
 
     function new (string name = "sys_scoreboard_1", uvm_component parent = null);
         super.new(name, parent);
     endfunction
 
 endclass