 class sys_scoreboard_5 extends uvm_component;
     `uvm_component_utils(sys_scoreboard_5)
 
     function new (string name = "sys_scoreboard_5", uvm_component parent = null);
         super.new(name, parent);
     endfunction
 
 endclass