package sys_scoreboard_pkg;

	import sys_seq_item_pkg::*;
	import uvm_pkg::*;
	`include "uvm_macros.svh"

	class sys_scoreboard extends uvm_scoreboard;
		`uvm_component_utils(sys_scoreboard)

		uvm_analysis_export #(sys_seq_item) sb_export;
		uvm_tlm_analysis_fifo #(sys_seq_item) sb_fifo;
		sys_seq_item seq_item_sb;
		
		int error_count=0;
		int correct_count=0;
		static int flag=0;
		static int counter=0;
		logic [7:0] frame;



			function new(string name="sys_scoreboard" , uvm_component parent=null);
				super.new(name,parent);
			endfunction

			function void build_phase(uvm_phase phase);
				super.build_phase(phase);
				sb_export=new("sb_export",this);
				sb_fifo=new("sb_fifo",this);

			endfunction

			function void connect_phase(uvm_phase phase);
				super.connect_phase(phase);
				sb_export.connect(sb_fifo.analysis_export);
			endfunction


			


			task run_phase(uvm_phase phase);
				super.run_phase(phase);
				forever begin
					sb_fifo.get(seq_item_sb);
				`uvm_info("score_board(sys_RX)",$sformatf("Done in sys DUT:%s",seq_item_sb.convert2string()),UVM_MEDIUM)
				end
			endtask

			function void report_phase(uvm_phase phase);
				super.report_phase(phase);
				`uvm_info("run_phase",$sformatf("totall successful transaction=%d",correct_count/2),UVM_MEDIUM)
				`uvm_info("run_phase",$sformatf("totall error transaction=%d",error_count/2),UVM_MEDIUM)
			endfunction

	endclass

endpackage 