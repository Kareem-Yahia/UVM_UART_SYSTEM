package global_pkg ;
		localparam EVEN=0;
		localparam ODD=1;
		localparam PAR_ENABLE=1;
		localparam PAR_DISABLE=0;
endpackage 