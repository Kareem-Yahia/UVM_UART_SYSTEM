package sys_sequence_pkg ;

	import sys_seq_item_pkg::*;
	import uvm_pkg::*;
	`include "uvm_macros.svh"

	class sys_sequence_reset extends uvm_sequence #(sys_seq_item);
		`uvm_object_utils (sys_sequence_reset)

		sys_seq_item seq_item;

		function new (string name="sys_sequence_reset");
			super.new(name);
		endfunction

		task body;
			seq_item = sys_seq_item::type_id::create ("seq_item");

			
			repeat(100) begin
				start_item (seq_item);
					assert(seq_item.randomize() with {seq_item.RST==0;seq_item.RX_IN==1;})
				finish_item(seq_item);
			end

		endtask

	endclass

	class sys_sequence_main extends uvm_sequence #(sys_seq_item);
		`uvm_object_utils (sys_sequence_main)

		sys_seq_item seq_item;

		function new (string name="sys_sequence_main");
			super.new(name);
		endfunction

		parameter EVEN=0;
		parameter ODD=1;
		parameter PAR_ENABLE=1;
		parameter PAR_DISABLE=0;
		bit parity_type;
		bit parity_enable;
		


		task body;
			seq_item = sys_seq_item::type_id::create ("seq_item");
			

			//////////////////////////////////////////////////////////////////////////////////////////////

			hold();
					Register_File_Write_command(2,8'b1000_01);
			hold();

			parity_type=EVEN;
			parity_enable=PAR_ENABLE;

			Register_File_Write_command(5,20,parity_type,parity_enable);
			Register_File_Write_command(6,25,parity_type,parity_enable);
			Register_File_Read_command(5,parity_type,parity_enable);
			Register_File_Read_command(6,parity_type,parity_enable);


			
			hold();
					Register_File_Write_command(2,8'b1000_11,parity_type,parity_enable);
			hold();
			parity_type=ODD;
			parity_enable=PAR_ENABLE;

			Register_File_Write_command(5,20,parity_type,parity_enable);
			Register_File_Write_command(6,25,parity_type,parity_enable);
			Register_File_Read_command(5,parity_type,parity_enable);
			Register_File_Read_command(6,parity_type,parity_enable);


			
			hold();
						Register_File_Write_command(2,8'b1000_00,parity_type,parity_enable);
			hold();
			parity_type=EVEN;
			parity_enable=PAR_DISABLE;

			Register_File_Write_command(5,20,parity_type,parity_enable);
			Register_File_Write_command(6,25,parity_type,parity_enable);
			Register_File_Read_command(5,parity_type,parity_enable);
			Register_File_Read_command(6,parity_type,parity_enable);



			///////////////////////////////////////////////////////////////////////////////////////////////
		endtask


		task send_specific_frame (input start,input [7:0] frame_t,input stop,input parity_type=EVEN,input parity_enable=1); // task used to send wrong frames
			  			uvm_resource_db#(logic [7:0])::set_override("*","frame_t", frame_t, this);

			 

			  start_item (seq_item);
				assert(seq_item.randomize() with {seq_item.RX_IN==start;seq_item.RST==1;})
			  finish_item(seq_item);

			for (int i = 0; i < 8; i++) begin
				 start_item (seq_item);
					assert(seq_item.randomize() with {seq_item.RX_IN==frame_t[i];seq_item.RST==1;})
			    finish_item(seq_item);
			end	

			if(parity_enable) begin
				if(parity_type==EVEN) begin
					start_item (seq_item);
						assert(seq_item.randomize() with {seq_item.RX_IN==^frame_t;seq_item.RST==1;})
			    	finish_item(seq_item);
				end
				else if(parity_type==ODD) begin
					start_item (seq_item);
						assert(seq_item.randomize() with {seq_item.RX_IN==~(^frame_t);seq_item.RST==1;})
			    	finish_item(seq_item);
				end
			end

			start_item (seq_item);
						assert(seq_item.randomize() with {seq_item.RX_IN==stop;seq_item.RST==1;})
			finish_item(seq_item);
		endtask

		task hold();
			start_item (seq_item);
						assert(seq_item.randomize() with {seq_item.RX_IN==1;seq_item.RST==1;})
			finish_item(seq_item);
		endtask



		task Register_File_Write_command (input [7:0] Address_t,input [7:0] DATA_t,input parity_type=EVEN,input parity_enable=1);

			send_specific_frame(0,'hAA,1,parity_type,parity_enable);
		
			send_specific_frame(0,Address_t,1,parity_type,parity_enable);

			send_specific_frame(0,DATA_t,1,parity_type,parity_enable);
		endtask

		task Register_File_Read_command (input [7:0] Address_t,input parity_type=EVEN,input parity_enable=1);
			
			send_specific_frame(0,'hBB,1,parity_type,parity_enable);
			
			send_specific_frame(0,Address_t,1,parity_type,parity_enable);

		endtask

		task ALU_Operation_command_with_operand (input [7:0] Operand_A_t,input [7:0] Operand_B_t,input [3:0] ALU_FUN_t,input parity_type=EVEN,input parity_enable=1);

			send_specific_frame(0,'hCC,1,parity_type,parity_enable);
			
			send_specific_frame(0,Operand_A_t,1,parity_type,parity_enable);
			
			send_specific_frame(0,Operand_B_t,1,parity_type,parity_enable);
			
			send_specific_frame(0,ALU_FUN_t,1,parity_type,parity_enable);
			
		endtask

		
		task ALU_Operation_command_with_No_operand (input [3:0] ALU_FUN_t,input parity_type=EVEN,input parity_enable=1);

		
			send_specific_frame(0,'hDD,1,parity_type,parity_enable);
			
			send_specific_frame(0,ALU_FUN_t,1,parity_type,parity_enable);

		endtask

	endclass

endpackage