package global_pkg ;
		localparam EVEN=0;
		localparam ODD=1;
		localparam PAR_ENABLE=1;
		localparam PAR_DISABLE=0;
		localparam PRESCALE_X8 = 8;
		localparam PRESCALE_X16 = 16;
		localparam PRESCALE_X32 = 32;

endpackage 